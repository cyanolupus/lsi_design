module test_vcs();
  initial begin
    $display("**************************");
    $display("****** Hello World! ******");
    $display("**************************");
    $finish;
  end
endmodule
